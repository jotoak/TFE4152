[aimspice]
[description]
2448
.include p18_model_card.inc
.include p18_cmos_models_tt.inc

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal
.param L1 = 0.36U
.param W1 = 5.04U
.param L2 = 1.08U
.param W2 = 1.08U
.param CC = 1.2pF
.param CS = 3pF

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1            ! Photo current source
d1 N1_R1C1 VDD dwell 1                        ! Reverse biased Diode
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40 ! Diode model
Cd1 N1_R1C1 VDD 30f                           ! Photo diode capacitor
.ends

xphoto 1 N1 Photodiode 
M1 N1 EXPOSE N2 0 NMOS L=L1 W=W1 
M2 N2 ERASE 0 0 NMOS L=L2 W=W2
M3 0 N2 N3 1 PMOS L=L1 W=W1
M4 N3 NRE_R1 OUT 1 PMOS L=L1 W=W1
CS N2 0 CS

xphoto2 1 N4 Photodiode 
M5 N4 EXPOSE N5 0 NMOS L=L1 W=W1 
M6 N5 ERASE 0 0 NMOS L=L2 W=W2
M7 0 N5 N6 1 PMOS L=L1 W=W1
M8 N6 NRE_R2 OUT 1 PMOS L=L1 W=W1
CS2 N5 0 CS

xphoto3 1 N7 Photodiode 
M9 N7 EXPOSE N8 0 NMOS L=L1 W=W1 
M10 N8 ERASE 0 0 NMOS L=L2 W=W2
M11 0 N8 N9 1 PMOS L=L1 W=W1
M12 N9 NRE_R1 OUT1 1 PMOS L=L1 W=W1
CS3 N8 0 CS

xphoto4 1 N10 Photodiode 
M13 N10 EXPOSE N11 0 NMOS L=L1 W=W1 
M14 N11 ERASE 0 0 NMOS L=L2 W=W2
M15 0 N11 N12 1 PMOS L=L1 W=W1
M16 N12 NRE_R2 OUT1 1 PMOS L=L1 W=W1
CS4 N11 0 CS

MC1 OUT OUT 1 1 PMOS L=L2 W=W2
CC1 OUT 0 CC

MC2 OUT1 OUT1 1 1 PMOS L=L2 W=W2
CC2 OUT1 0 CC



.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(OUT1) V(OUT)







[tran]
0.1
60ms
X
X
0
[ana]
4 0
[end]
